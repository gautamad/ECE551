module Mul();

wire signed [14:0] a,b;
wire signed [29:0] c;

assign c = a * b;

endmodule
