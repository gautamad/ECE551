module ALU_tb();
	
	reg 

endmodule
