library verilog;
use verilog.vl_types.all;
entity add4bit_tb is
end add4bit_tb;
