library verilog;
use verilog.vl_types.all;
entity Mul is
end Mul;
