library verilog;
use verilog.vl_types.all;
entity osc_tb is
end osc_tb;
