library verilog;
use verilog.vl_types.all;
entity PWM_tb is
end PWM_tb;
