library verilog;
use verilog.vl_types.all;
entity add8bit_tb is
end add8bit_tb;
