library verilog;
use verilog.vl_types.all;
entity osc is
    port(
        en              : in     vl_logic;
        \out\           : out    vl_logic
    );
end osc;
