module A2D_intf();

endmodule