library verilog;
use verilog.vl_types.all;
entity moto_driver_tb is
end moto_driver_tb;
