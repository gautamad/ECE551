library verilog;
use verilog.vl_types.all;
entity BarCode_tb is
end BarCode_tb;
