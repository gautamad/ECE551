library verilog;
use verilog.vl_types.all;
entity UART_rx_tb is
end UART_rx_tb;
